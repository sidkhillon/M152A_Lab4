module Countdown(
    input wire clk,
    input wire clk_countdown,
    input wire rst,
    input wire start,
    output reg [1:0] anode,
    output reg countdown_done,
    output reg countdown_in_action
);

reg start_sync1, start_sync2;  
reg start_pulse;

always @(posedge clk_countdown or posedge rst) begin
    if (rst) begin
        start_sync1 <= 0;
        start_sync2 <= 0;
    end else begin
        start_sync1 <= start;
        start_sync2 <= start_sync1;
    end
end

always @(posedge clk_countdown or posedge rst) begin
    if (rst)
        start_pulse <= 0;
    else
        start_pulse <= start_sync2 & ~start_pulse;
end

always @(posedge clk_countdown or posedge rst) begin
    if (rst) begin
        anode <= 2'b00;
        countdown_done <= 0;
        countdown_in_action <= 0;
    end else if (start_pulse) begin
        anode <= 2'b00;
        countdown_done <= 0;
        countdown_in_action <= 1;
    end else if (countdown_in_action) begin
        if (anode == 2'd3) begin
            countdown_done <= 1;
            countdown_in_action <= 0;
        end else begin
            anode <= anode + 1;
            countdown_done <= 0;
        end
    end else begin
        countdown_done <= 0;
    end
end

endmodule
